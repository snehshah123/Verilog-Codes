// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Thu Mar 28 07:09:48 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module sneh91 (
    CLK,RST,X,
    Z);

    input CLK;
    input RST;
    input X;
    tri0 RST;
    tri0 X;
    output Z;
    reg Z;
    reg reg_Z;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter S0=0,S1=1,S2=2,S3=3;

    initial
    begin
        reg_Z <= 1'b0;
    end

    always @(posedge CLK)
    begin
        if (CLK) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or RST or X or reg_Z)
    begin
        if (RST) begin
            reg_fstate <= S0;
            reg_Z <= 1'b0;
            Z <= 1'b0;
        end
        else begin
            reg_Z <= 1'b0;
            Z <= 1'b0;
            case (fstate)
                S0: begin
                    if ((X == 1'b1))
                        reg_fstate <= S1;
                    else if ((X == 1'b0))
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;
                end
                S1: begin
                    if ((X == 1'b0))
                        reg_fstate <= S2;
                    else if ((X == 1'b1))
                        reg_fstate <= S1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S1;
                end
                S2: begin
                    if ((X == 1'b0))
                        reg_fstate <= S0;
                    else if ((X == 1'b1))
                        reg_fstate <= S3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S2;
                end
                S3: begin
                    if ((X == 1'b1))
                        reg_fstate <= S1;
                    else if ((X == 1'b0))
                        reg_fstate <= S2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S3;

                    if ((X == 1'b1))
                        reg_Z <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_Z <= 1'b0;
                end
                default: begin
                    reg_Z <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
            Z <= reg_Z;
        end
    end
endmodule // sneh91
